// module websocket
