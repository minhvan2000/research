// module main

// import time
// import log

// // Setup Logger
// fn (mut app App) setup_logger() {
// 	handle.logger.set_level(.debug)

// 	handle.logger.set_full_logpath('./src/logs/log_${time.now().ymmdd()}.log')
// 	handle.logger.log_to_console_too()
// }

// pub fn (mut app App) warn(msg string) {
// 	handle.logger.warn(msg)

// 	handle.logger.flush()
// }

// pub fn (mut app App) info(msg string) {
// 	handle.logger.info(msg)

// 	handle.logger.flush()
// }

// pub fn (mut app App) debug(msg string) {
// 	handle.logger.debug(msg)

// 	handle.logger.flush()
// }
